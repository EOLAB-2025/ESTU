parameter SPIKE_MEM_WIDTH      = 4;
parameter SPIKE_MEM_DEPTH      = 1024;
parameter RAM_PERFORMANCE      = "HIGH_PERFORMANCE";
parameter INIT_FILE_SM1        = "C:/Users/Mauro/Desktop/Mauro/Borsa/Spikeformer/Spikeformer/scripts/INIT_FILE_SM1.txt";
parameter INIT_FILE_SM2        = "C:/Users/Mauro/Desktop/Mauro/Borsa/Spikeformer/Spikeformer/scripts/INIT_FILE_SM2.txt";
parameter INIT_FILE_SM3        = "C:/Users/Mauro/Desktop/Mauro/Borsa/Spikeformer/Spikeformer/scripts/INIT_FILE_SM3.txt";
parameter INIT_FILE_SM4        = "C:/Users/Mauro/Desktop/Mauro/Borsa/Spikeformer/Spikeformer/scripts/INIT_FILE_SM4.txt";
parameter NUM_MEMS_SPIKE_MEM   = 4;
parameter DEPTH_INT_MEM        = 1024;
parameter INIT_FILE_INTMEM1    = "C:/Users/Mauro/Desktop/Mauro/Borsa/Spikeformer/Spikeformer/scripts/INIT_FILE_INTMEM1.txt";
parameter INIT_FILE_INTMEM2    = "C:/Users/Mauro/Desktop/Mauro/Borsa/Spikeformer/Spikeformer/scripts/INIT_FILE_INTMEM2.txt";
parameter DIM_ADDR_SPIKE_MEM   = 12;
parameter DIM_ADDR_SPRAM       = 14;
parameter DIM_MAX_MEM          = 14;
parameter DIM_INPUT_NEURONS    = 5;
parameter DIM_OUTPUT_NEURONS   = 10;
parameter DIM_MAX_LOGIC_ADDRESS= 10;
parameter DEPTH_STACK          = 3468;
parameter INIT_STACK           = "C:/Users/Mauro/Desktop/Mauro/Borsa/Spikeformer/Spikeformer/scripts/stack_init.txt";
parameter DATA_WIDTH           = 8;
parameter V_COMP_K_Q           = 800;
parameter WIDTH_BRAM           = 4;
parameter WIDTH_SPRAM          = 16;
parameter DIM_MODE             = 5;
parameter DIM_GROUP_SPIKES     = 2;
parameter DIM_SUMS_SPIKES      = 16;
parameter NUM_MEMS             = 4;
parameter DIM_OFFSET           = 6;
parameter DIM_GROUP_SPIKE4     = 4;
parameter DIM_GROUP_16         = 16;
parameter DIM_CURRENT          = 22;
parameter DIM_CTRL             = 7;
parameter NEURON               = 256;
parameter DIM_CURR_DECAY_LIF   = 14;
parameter DIM_VOLT_DECAY_LIF   = 14;
parameter WIDTH_LIF            = 23;
parameter INSTR_MEM_WIDTH      = 32;
parameter TOT_NUM_INSTR        = 30;
parameter DIM_INSTR            = 179;
parameter NUM_INSTR            = 6;
parameter DIM_NUM_INSTR        = 3;
parameter INSTR_MEM_DEPTH      = 180;
parameter INIT_INSTR_MEM       = "C:/Users/Mauro/Desktop/Mauro/Borsa/Spikeformer/Spikeformer/scripts/instr_mem.txt";

