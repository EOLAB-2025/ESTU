`timescale 1ns / 1ps

module wr_controller #(
    parameter DATA_WIDTH = 8,   // Data width
    parameter P_SPRAM = 2, // Number of parallel data
    parameter P_BRAM = 2, // Number of parallel group of spikes
    parameter DIM_MODE = 4,
    parameter WIDTH_BRAM = 4,
    parameter WIDTH_SPRAM = 16,
    parameter DIM_TIMESTEP = 8
)(
    // External signals
    // input [3:0] ext_ctrl,
    // input [WIDTH_SPRAM-1:0] ext_datain_spram1,
    // input [WIDTH_SPRAM-1:0] ext_datain_spram2,
    // input [WIDTH_BRAM-1:0] ext_datain_bram1,
    // input [WIDTH_BRAM-1:0] ext_datain_bram2,
    // Accelerator signals
    input clk,
    input rst,
    input clr,
    input en, // Enable signal
    input valid_data, // Valid data signal
    input [DATA_WIDTH-1:0] data_int, // Integer data of 8 bit width. Output of the matmul(spike,spike) operation
    input [DATA_WIDTH*2-1:0] sum_spikes,
    input [1:0] spike_out, // Output of the LIF neuron
    input [DIM_MODE-1:0] mode, // Mode of the operation
    input [DIM_TIMESTEP-1:0] timestep,
    input [3:0] group_in_spikes,
    input new_spike,  // 1 bit signal that represents the new spike generated by the LIF neuron
    input use_v,
    input v_gen_id,
    input [1:0] sel_data_int, // Forse da togliere
    input clr_valid_ll_ext, // Clear valid last layer output
    input last_layer, 
    input valid_instr,
    output wren_bram1, // Write enable signal for the BRAM 1
    output wren_bram2, // Write enable signal for the BRAM 2
    output wren_spram1, // Write enable signal for the SPRAM 1
    output wren_spram2, // Write enable signal for the SPRAM 2
    output [WIDTH_BRAM - 1 : 0] data_in_bram1,
    output [WIDTH_BRAM - 1 : 0] data_in_bram2,
    output [WIDTH_SPRAM - 1 : 0] data_in_spram1,
    output [WIDTH_SPRAM - 1 : 0] data_in_spram2,
    output active_group_out,
    output matmul_ss,
    output valid_last_layer_output,
    output [12:0] output_last_layer

);
    // Internal signals
    wire [3:0] data_out_V;
    wire sel_mux_V [3:0];
    wire [DATA_WIDTH - 1 : 0] data_out_int [3:0];
    `ifdef SIMULATION
    wire [DATA_WIDTH-1 : 0] data_out_intsim1;
    wire [DATA_WIDTH-1 : 0] data_out_intsim2;
    wire [DATA_WIDTH-1 : 0] data_out_intsim3;
    wire [DATA_WIDTH-1 : 0] data_out_intsim4;
    assign data_out_intsim1 = data_int_reg[0];
    assign data_out_intsim2 = data_int_reg[1];
    assign data_out_intsim3 = data_int_reg[2];
    assign data_out_intsim4 = data_int_reg[3];
    `endif
    // ---------------------------- S2P Int writing --------------------------------------
    // Used only for matmul(spike,spike) operation
    // -------------------------------------------------------------------------
    assign matmul_ss = ~(|mode)&en;
    reg [DATA_WIDTH-1:0] data_int_reg [3:0];
    always @(posedge clk) begin
        if (rst | clr) begin
            data_int_reg[0] <= 0;
            data_int_reg[1] <= 0;
            data_int_reg[2] <= 0;
            data_int_reg[3] <= 0;
        end 
        else if (valid_data) begin
            data_int_reg[0] <= data_out_int[0];
            data_int_reg[1] <= data_out_int[1];
            data_int_reg[2] <= data_out_int[2];
            data_int_reg[3] <= data_out_int[3];
        end
    end
    wire sel_data_int_mux [3:0];
    
    assign sel_data_int_mux[0] = ~sel_data_int[1] &  ~sel_data_int[0];
    assign sel_data_int_mux[1] = ~sel_data_int[1] &  sel_data_int[0];
    assign sel_data_int_mux[2] = sel_data_int[1] &  ~sel_data_int[0];
    assign sel_data_int_mux[3] = sel_data_int[1] &  sel_data_int[0];

    assign data_out_int[0] = sel_data_int_mux[0] ? data_int : data_int_reg[0];
    assign data_out_int[1] = sel_data_int_mux[0] ? 8'b0 : (sel_data_int_mux[1] ? data_int : data_int_reg[1]);
    assign data_out_int[2] = sel_data_int_mux[0] ? 8'b0 : (sel_data_int_mux[2] ? data_int : data_int_reg[2]);
    assign data_out_int[3] = sel_data_int_mux[0] ? 8'b0 : (sel_data_int_mux[3] ? data_int : data_int_reg[3]);
    // ---------------------------- End S2P Int writing --------------------------------------
    
    // ---------------------------- S2P Spikes writing --------------------------------------
    wire [2*P_BRAM-1:0] data_out_s2p_bram;
    wire valid_s2p_bram;
    s2p_rev #(
        .P(P_BRAM),
        .DATA_IN(2)
    ) s2p_instance_bram (
        .clk(clk),
        .rst(rst | clr),
        .en(valid_data & mode[3]),
        .data_in(spike_out),
        .data_out(data_out_s2p_bram),
        .valid(valid_s2p_bram)
    ); 
    // ---------------------------- End S2P Spikes writing --------------------------------------

    // ---------------------------- Write of V --------------------------------------
    assign sel_mux_V[0] = ~timestep[0] &  ~timestep[1];
    assign sel_mux_V[1] = timestep[0] &  ~timestep[1];
    assign sel_mux_V[2] = ~timestep[0] &  timestep[1];
    assign sel_mux_V[3] = timestep[0] &  timestep[1];

    assign data_out_V[0] = sel_mux_V[0] ? 1'b0 : (sel_mux_V[3] ? new_spike : group_in_spikes[0]);
    assign data_out_V[1] = sel_mux_V[0] ? 1'b0 : (sel_mux_V[2] ? new_spike : group_in_spikes[1]);
    assign data_out_V[2] = sel_mux_V[0] ? 1'b0 : (sel_mux_V[1] ? new_spike : group_in_spikes[2]);
    assign data_out_V[3] = sel_mux_V[0] ? new_spike : group_in_spikes[3];
    
    wire ored_spikes;
    assign ored_spikes = |group_in_spikes;
    wire ored_data_in_bram = |data_in_bram1;
    assign active_group_out = v_gen_id ? (sel_mux_V[0] ? new_spike : (ored_spikes ? 1'b0 : new_spike)) : (ored_data_in_bram & ~v_gen_id);
    // ---------------------------- End Write of V --------------------------------------

    // ---------------------------- Last Layer -----------------------------------------

    reg [12:0] ctrl_reg_ll;
    wire clr_ll;
    assign clr_ll = (valid_instr & last_layer);
    reg [12:0] dout_ll;
    reg valid_dout_ll;
    wire en_last_layer;
    assign en_last_layer = valid_data & last_layer & ~clr_ll;
    always @(posedge clk) begin
        if (rst)
            ctrl_reg_ll <= 0;
        else if (clr_ll | clr_valid_ll_ext)
            ctrl_reg_ll <= 1;
        else if (en_last_layer)
            ctrl_reg_ll <= ctrl_reg_ll<<1;
    end
    integer i;
    always @(posedge clk) begin
        if (rst | clr_ll )
            dout_ll <= 0;
        else if (en_last_layer)
            for (i=0; i<13; i=i+1) begin
                if (ctrl_reg_ll[i])
                    dout_ll[i] <= new_spike;
                else
                    dout_ll[i] <= dout_ll[i];
            end
    end

    always @(posedge clk) begin
        if (rst | clr_ll)
            valid_dout_ll <= 0;
        else 
            valid_dout_ll <= ctrl_reg_ll[12]&en_last_layer;
    end

    assign output_last_layer = dout_ll;
    assign valid_last_layer_output = valid_dout_ll;
    // ---------------------------- End Last Layer -----------------------------------------

    // Output assignments
    assign wren_bram1 = v_gen_id ?  valid_data : valid_s2p_bram;
    assign wren_bram2 = v_gen_id ? valid_data : valid_s2p_bram;
    assign wren_spram1 = valid_data;
    assign wren_spram2 = valid_data;
    
    // MUX DATA IN
    assign data_in_bram1 = ((v_gen_id) ? data_out_V : data_out_s2p_bram);
    assign data_in_bram2 = ((v_gen_id) ? data_out_V : data_out_s2p_bram);
    assign data_in_spram1 =  ({mode[2]} ? sum_spikes : {data_out_int[0],data_out_int[1]});
    assign data_in_spram2 = ({mode[2]} ? sum_spikes : {data_out_int[2],data_out_int[3]});
    
    ////////////////////////////
    //  _               ____  //
    // | | ___   __ _  |___ \ //
    // | |/ _ \ / _` |   __)  //
    // | | (_) | (_| |  / __/ //
    // |_|\___/ \__, | |_____ //
    //          |___/         //
    ////////////////////////////
    
    //  The following function calculates the address width based on specified RAM depth
    function integer clogb2;
    input integer depth;
        for (clogb2=0; depth>0; clogb2=clogb2+1)
        depth = depth >> 1;
    endfunction 
endmodule