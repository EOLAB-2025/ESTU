`timescale 1ns / 1ps


module datapath #(
    parameter DIM_MODE = 5,
    parameter DIM_GROUP_SPIKE4 = 4, // Most of the operations such as dense(spike,int) are done in groups of 4
    parameter DIM_GROUP_16 = 16, // matmul(spike,spike) is done in groups of 16
    parameter DATA_WIDTH = 8, // Data width of int data
    parameter NUM_MEMS = 4,
    parameter DIM_CURRENT = 22,
    parameter DIM_CTRL = 7,
    // LIF Section
    parameter NEURON = 717,
    parameter DIM_CURR_DECAY_LIF = 14,
    parameter DIM_VOLT_DECAY_LIF = 14,
    parameter WIDTH_LIF = 23
)(
    input clk, rst, valid_inference, acc_clear_and_go, block_rd_cnt_lif, clr, en,
    input [DIM_CTRL - 1 : 0] ctrl_sig, 
    input use_v, empty,
    input [DIM_MODE - 1 : 0] mode,
    input [DIM_GROUP_SPIKE4 - 1 : 0] spikes_in_1, spikes_in_2, // Group of 4 spikes used for dense(spike,int), sum(spike,spike) and sum(spike,int)
    input [DIM_GROUP_16 - 1 : 0] spikes_in16_1, spikes_in16_2, // Groups of 16 spikes used for matmul(spike,spike)
    input [DIM_GROUP_16 - 1 : 0] data_int1, data_int2, // 2 Groups of 2 8 bit integers, output of the int mem
    input [NUM_MEMS-1 : 0] r_en_mems,
    input [DIM_VOLT_DECAY_LIF - 1 : 0] voltage_decay,
    input [WIDTH_LIF - 1 : 0] threshold,
    input use_stack,
    input v_gen_id,
    input valid_op_mmu,
    input last_layer,
    output spike_s_out, // One bit signal that represents the new spike generated by the LIF neuron. Used for the V generation writing phase
    output [1:0] spike_p_out, // Output of the LIF neuron. Used in all the dense operations except for the V generation writing phase
    output [DATA_WIDTH - 1 : 0] data_int_out,
    output [DATA_WIDTH*2 - 1 : 0] data_int_out_sums,
    output valid_datapath,
    output valid_int_neuron // Valid signal for the LIF neuron output
);

    // Local parameters
    localparam SUM = DIM_GROUP_SPIKE4/2;
    localparam DIM_POP_CNT = clogb2(DIM_GROUP_16);
    // Groups of 4 spikes 
    wire [DATA_WIDTH-1:0] spike_a1 [SUM-1:0]; 
    wire [DATA_WIDTH-1:0] spike_b1 [SUM-1:0];   
    wire [DATA_WIDTH-1:0] spike_a2 [SUM-1:0]; 
    wire [DATA_WIDTH-1:0] spike_b2 [SUM-1:0];  
    // Groups of 2 data int of 8 bits
    wire signed [DATA_WIDTH-1:0] weights_a [SUM-1:0]; 
    wire signed [DATA_WIDTH-1:0] weights_b [SUM-1:0]; 
    // 4 MUX pre AND for spikes selection
    wire [DATA_WIDTH - 1: 0] mux_out_spike_b [SUM-1:0];
    wire [DATA_WIDTH - 1: 0] mux_out_spike_a [SUM-1:0]; 
    wire [DATA_WIDTH - 1: 0] mux_out_spike_b2 [SUM-1:0];
    wire [DATA_WIDTH - 1: 0] mux_out_spike_a2 [SUM-1:0]; 
    // 4 8 bit ANDs: used for dense(spike,int) operation
    wire [DATA_WIDTH - 1 : 0] and_out_b [SUM-1:0];
    wire [DATA_WIDTH - 1 : 0] and_out_a [SUM-1:0];
    //4 MUX used to control the routing for sum(spike,spike) and sum(spike,int) operations
    wire [DATA_WIDTH - 1: 0] mux_out_sum_1 [SUM-1:0];
    reg [DATA_WIDTH - 1: 0] mux_out_sum_2 [SUM-1:0];
    // 4 MUX for the selection of the Accumulator input
    wire [DATA_WIDTH - 1: 0] mux_out_acc_a [SUM-1:0];
    wire [DATA_WIDTH - 1: 0] mux_out_acc_b [SUM-1:0];
    // Adder SIMD: perform the pairwise addition
    wire signed [DATA_WIDTH:0] double_adder_out [SUM-1:0]; // Forse da cambiare la dimensione
    wire double_adder_en;
    // Accumulator
    wire signed [WIDTH_LIF-1:0] acc_out;
    wire signed [WIDTH_LIF-2:0] acc_in [SUM-1:0];
    wire c_en_acc [2:0]; // NOTA: FARE L'ASSIGN OPPORTUNAMENTE DA CTRL_SIG!!!!!!!!!
    // Multipliers
    wire signed [2*DATA_WIDTH-1 : 0] prod_a, prod_b;
    reg signed [2*DATA_WIDTH-1 : 0] prod_a_r, prod_b_r;
    // Matmul spike spike
    reg [DIM_POP_CNT-1:0] pop_cnt_r;
    wire [DIM_POP_CNT-1:0] pop_cnt;
    wire [DIM_GROUP_16 - 1 : 0] and_16;
    // Other control signals
    reg en_d;
    // LIF Unit
    localparam WEIGHT = 8; 
    wire valid_neuron;
    wire en_neuron;
    wire en_lif; // Fare l'assign in base al ctrl_sig
    reg en_neuron_d;
    wire [WIDTH_LIF - 1 : 0] neuron_lp_voltage;
    // For generate statement
    genvar i;



    // Spike sorting group 1
    generate
    for (i = 0; i < SUM; i = i + 1) begin 
        assign spike_a1[i] = empty ? {DATA_WIDTH{1'b0}} : {(DATA_WIDTH){spikes_in_1[i + SUM]}};
        assign spike_b1[i] = empty ? {DATA_WIDTH{1'b0}} : {(DATA_WIDTH){spikes_in_1[i]}};
    end
    endgenerate

    // Spike sorting group 2   
    generate
        for (i = 0; i < SUM; i = i + 1) begin 
            assign spike_a2[i] = empty ? {DATA_WIDTH{1'b0}} : {(DATA_WIDTH){spikes_in_2[i + SUM]}};
            assign spike_b2[i] = empty ? {DATA_WIDTH{1'b0}} : {(DATA_WIDTH){spikes_in_2[i]}};
        end
    endgenerate

    // Data int sorting 
    generate
        for (i = 0; i < SUM; i = i + 1) begin 
            assign weights_a[i] = data_int1[(i+1)*DATA_WIDTH-1 -: DATA_WIDTH];       
            assign weights_b[i] = data_int2[(i+1)*DATA_WIDTH-1 -: DATA_WIDTH];       
        end
    endgenerate

    `ifdef SIMULATION
        wire [DATA_WIDTH - 1: 0] weight_sim1a, weight_sim1b, weight_sim2a, weight_sim2b;
        wire [DATA_WIDTH-1:0] and_out_sim1a, and_out_sim1b, and_out_sim2a, and_out_sim2b;
        assign and_out_sim1a = and_out_a[0];
        assign and_out_sim1b = and_out_b[0];
        assign and_out_sim2a = and_out_a[1];
        assign and_out_sim2b = and_out_b[1];
        assign weight_sim1a = weights_a[0];
        assign weight_sim1b = weights_b[0];
        assign weight_sim2a = weights_a[1];
        assign weight_sim2b = weights_b[1];
    `endif


    // 4 MUX pre AND for spikes selection
    assign mux_out_spike_b[0] = r_en_mems[1] ? spike_b2[0] : spike_b1[0];
    assign mux_out_spike_b[1] = r_en_mems[1] ? spike_b2[1] : spike_b1[1];
    assign mux_out_spike_a[0] = r_en_mems[1] ? spike_a2[0] : spike_a1[0];
    assign mux_out_spike_a[1] = r_en_mems[1] ? spike_a2[1] : spike_a1[1];


    // 4 8 bit ANDs: used for dense(spike,int) operation
    assign  and_out_b[0] = mux_out_spike_b[0] & weights_b[0];
    assign  and_out_b[1] = mux_out_spike_b[1] & weights_b[1];
    assign  and_out_a[0] = mux_out_spike_a[0] & weights_a[0];
    assign  and_out_a[1] = mux_out_spike_a[1] & weights_a[1];

    //4 MUX used to control the routing for sum(spike,spike) and sum(spike,int) operations
    // Pairwise selection in groups of odd/even indices
    /*
    assign mux_out_sum_1[0] = en ? {7'b0, spike_b1[1][0]} : {7'b0, spike_b1[0][0]};
    assign mux_out_sum_1[1] = en ? {7'b0, spike_a1[1][0]} : {7'b0, spike_a1[0][0]};
    always @(*) begin
        case ({mode[4], en})
            2'b00: begin
                mux_out_sum_2[0] = {7'b0, spike_b2[0][0]};
                mux_out_sum_2[1] = {7'b0, spike_a2[0][0]};
            end
            2'b01: begin
                mux_out_sum_2[0] = {7'b0, spike_b2[1][0]};
                mux_out_sum_2[1] = {7'b0, spike_a2[1][0]};
            end
            2'b10: begin
                mux_out_sum_2[0] = weights_b[0];
                mux_out_sum_2[1] = weights_a[0];
            end
            2'b11: begin
                mux_out_sum_2[0] = weights_b[1];
                mux_out_sum_2[1] = weights_a[1];
            end
        endcase    
    end
    */
    assign mux_out_sum_1[0] = en ?  {7'b0, spike_a1[0][0]} : {7'b0, spike_b1[0][0]};
    assign mux_out_sum_1[1] = en ?  {7'b0, spike_a1[1][0]} : {7'b0, spike_b1[1][0]};

    wire [7:0] mux_out_sum_weigths [1:0];

    assign mux_out_sum_weigths[0] = r_en_mems[2] ? weights_a[0] : weights_b[0];
    assign mux_out_sum_weigths[1] = r_en_mems[2] ? weights_a[1] : weights_b[1];

    always @(*) begin
        case ({mode[4], en})
            2'b00: begin
                mux_out_sum_2[0] = {7'b0, spike_b2[0][0]};
                mux_out_sum_2[1] = {7'b0, spike_b2[1][0]};
            end
            2'b01: begin
                mux_out_sum_2[0] = {7'b0, spike_a2[0][0]};
                mux_out_sum_2[1] = {7'b0, spike_a2[1][0]};
            end
            2'b10: begin
                mux_out_sum_2[0] = mux_out_sum_weigths[0];
                mux_out_sum_2[1] = mux_out_sum_weigths[1];
            end
            2'b11: begin
                mux_out_sum_2[0] = mux_out_sum_weigths[0];
                mux_out_sum_2[1] = mux_out_sum_weigths[1];
            end
        endcase    
    end

    // 4 MUX for the selection of the Accumulator input
    assign mux_out_acc_a[0] = mode[2] ? mux_out_sum_1[0] : and_out_a[0];
    assign mux_out_acc_a[1] = mode[2] ? mux_out_sum_1[1] : and_out_a[1];
    assign mux_out_acc_b[0] = mode[2] ? mux_out_sum_2[0] : and_out_b[0];
    assign mux_out_acc_b[1] = mode[2] ? mux_out_sum_2[1] : and_out_b[1];

    // Control for the sum operations
    // Delayed enable
    always @(posedge clk) begin
        if (rst | clr) 
            en_d <= 0;
        else
            en_d <= en;
    end

    // Adder SIMD: perform the pairwise addition 
    assign double_adder_en = en_d&(mode[2]) | en;
    adder_simd #(SUM, DATA_WIDTH)
        double_adder_inst
        (
        clk,
        double_adder_en,
        clr,
        mux_out_acc_a[0],
        mux_out_acc_a[1],
        mux_out_acc_b[0],
        mux_out_acc_b[1],
        double_adder_out[0],
        double_adder_out[1]
    );

    // Accumulator: used for all the dense operations and for the matmul(spike,int) operation
    // Mux accumulator: used to select the input of the accumulator -> it can be the output of the double adder or the output of the multiplier
    assign acc_in[0] = mode[0] ? prod_a_r : double_adder_out[0];
    assign acc_in[1] = mode[0] ? prod_b_r : double_adder_out[1];
    assign c_en_acc[0] = use_stack ? (use_v ? ctrl_sig[3]|ctrl_sig[4] : ctrl_sig[5]) : ctrl_sig[2];
    assign c_en_acc[1] = use_stack ? (use_v ? ctrl_sig[4]|ctrl_sig[5] : ctrl_sig[6]) : ctrl_sig[3];
    assign c_en_acc[2] = use_stack ? (use_v ? ctrl_sig[5]|ctrl_sig[6] : ctrl_sig[7]) : ctrl_sig[4];
    accumulator
    #(WIDTH_LIF-1)
    accumulator_inst
    (
    clk,c_en_acc[0],c_en_acc[1],c_en_acc[2],(rst),(use_v ? 1'b0: acc_clear_and_go),(use_v ? (acc_clear_and_go|clr) : clr),acc_in[0],acc_in[1],acc_out
    );

    // Multipliers
    assign prod_a = weights_a[0] * weights_b[0];
    assign prod_b = weights_a[1] * weights_b[1];
    always @(posedge clk) begin
        if (rst | clr) begin
            prod_a_r <= 0;
            prod_b_r <= 0;
        end
        else begin
            prod_a_r <= prod_a;
            prod_b_r <= prod_b;
        end
    end

    // 16 ANDs: This section is used only for the matmul(spike,spike) operation
    generate 
        for (i = 0; i < 16; i = i + 1) begin : ands
            assign and_16[i] = spikes_in16_1[i] & spikes_in16_2[i];
        end
    endgenerate
    // Population counter
    assign pop_cnt = and_16[0] + and_16[1] + and_16[2] + and_16[3] + and_16[4] + and_16[5] + and_16[6] + and_16[7] + and_16[8] + and_16[9] + and_16[10] + and_16[11] + and_16[12] + and_16[13] + and_16[14] + and_16[15];
    always @(posedge clk) begin
        if (rst | clr) begin
            pop_cnt_r <= 0;
        end
        else begin
            pop_cnt_r <= pop_cnt;
        end
    end


    // -------------------------------------------- LIF MODULE --------------------------------------------
    always @(posedge clk) begin
        if (rst | clr) begin
            en_neuron_d <= 0;
        end
        else begin
            en_neuron_d <= en_neuron;
        end
    end
    assign en_lif = acc_clear_and_go;
    assign en_neuron = en_lif & mode[3] & ~valid_op_mmu;
    neuron_lp 
    #(.DEPTH(NEURON),.WIDTH(WIDTH_LIF),.WEIGHT(WEIGHT))
     neuron_lp_i
        (
        .clk(clk), 
        .rst(rst | clr),
        .rst_fifo(valid_inference |  rst), 
        .en(en_neuron), 
        .en_d(en_neuron_d),
        .voltage_decay(voltage_decay), .threshold(threshold), 
        .block_rd_cnt_lif(block_rd_cnt_lif),
        .synaptic_current(acc_out),
        .valid(valid_neuron),
        .spike_p(spike_p_out),
        .voltage_ready(valid_int_neuron),
        .voltage(neuron_lp_voltage),
        .spike_s(spike_s_out)
        );

    // Output assignments
    assign data_int_out = pop_cnt_r; 
    assign data_int_out_sums = {double_adder_out[1][DATA_WIDTH-1 -: DATA_WIDTH], double_adder_out[0][DATA_WIDTH-1 -: DATA_WIDTH]};
    assign valid_datapath = (v_gen_id|last_layer) ? valid_int_neuron : valid_neuron;

    ////////////////////////////
    //  _               ____  //
    // | | ___   __ _  |___ \ //
    // | |/ _ \ / _` |   __)  //
    // | | (_) | (_| |  / __/ //
    // |_|\___/ \__, | |_____ //
    //          |___/         //
    ////////////////////////////
    
    //  The following function calculates the address width based on specified RAM depth
    function integer clogb2;
    input integer depth;
        for (clogb2=0; depth>0; clogb2=clogb2+1)
        depth = depth >> 1;
    endfunction  
endmodule